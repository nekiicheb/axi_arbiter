`include "globals.vh"

interface AxiAddition (
  input logic aclk

);
	logic [`CHANNELS_W-1:0] idx_channel
/* modport In(input aclk );
modport Out(input aclk, input areset_n); */

endinterface