`ifndef GLOBALS
`define GLOBALS

/* `define DATA_SIZE  32
`define ID_SIZE    8
`define CHANNELS_W 2
`define NUM_CHANNELS 4
`define MAX_PACKET_SIZE 4 */

`endif
